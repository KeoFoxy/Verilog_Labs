module lab_3_individual (sw, hex0, hex1, hex2, hex3, x ,y);
input [4:0] sw;

output reg [6:0] hex0;
output reg [6:0] hex1;
output [6:0] hex2;
output [6:0] hex3;
output reg [6:0] x; //переменная для хранения десятичных значений
output reg [6:0] y; //все числа от 0 -> 9

//Сделаем по красоте и остальные неиспользованные 
//индикаторы как 0 0
assign hex3 = 7'b1000000;
assign hex2 = 7'b1000000;


always @*
begin

    //Далее хреначим числа
    //Обозначим, с каким числом работаем
    //С 10 20 30 или 0-9

    if(sw[4:0] > 29)
    x = 3;
    else if(sw[4:0] > 19)
    x = 2;
    else if(sw[4:0] > 9)
    x = 1;
    else 
    x = 0;

    //Выводим число, отвечающее за десятки
    case(x)
    0:hex1 =7'b1000000;
    1:hex1 =7'b1001111;
    2:hex1 =7'b0100100;
    3:hex1 =7'b0110000;
    endcase
    //Далее выкидаем из числа 10ки и получаем число от 0->9
    //
    y = sw[4:0]-x*10;

    //Далее передаем в кейс и он уже нарисует нам число, 
    //аналогично прошлым задания в лабе
    case(y)
    0:hex0=7'b1000000;
    1:hex0=7'b1001111;
    2:hex0=7'b0100100;
    3:hex0=7'b0110000;
    4:hex0=7'b0011001;
    5:hex0=7'b0010010;
    6:hex0=7'b0000010;
    7:hex0=7'b1111000;
    8:hex0=7'b0000000;
    9:hex0=7'b0010000;
    endcase
end

endmodule