module lab_3_3_1 (sw, ledg);
input [7:0] sw;
output reg [7:0] ledg;

//сначала забираем десятку у числа
//Смотрим какое число формируют свичи в битках
//от 1 до 9
//Далее мы берем и по прнципу работы BTD добикидываем к ним числа от 0-9
//чтобы сформировать двузначное число
//Далее
//Для примера
//69 = вы снимаем первых четрых свитчей 6, далее по кейсу
//мы закинем 9ку
//Верилог умный, он сам там все преобразует

always @*
begin
case (sw[7:4])
    0:ledg= 0+sw[3:0];
    1:ledg=10+sw[3:0];
    2:ledg=20+sw[3:0];
    3:ledg=30+sw[3:0];
    4:ledg=40+sw[3:0];
    5:ledg=50+sw[3:0];
    6:ledg=60+sw[3:0];
    7:ledg=70+sw[3:0];
    8:ledg=80+sw[3:0];
    9:ledg=90+sw[3:0];
endcase
end                                                           

endmodule  