module lab_3_3_1 (sw, ledg);
input [7:0] sw;
output [7:0] ledg;

wire [7:0] dozens = sw[7:4];
wire [3:0] ones = sw[3:0];

reg [7:0] temp;

always @*
begin
case (sw[7:4])
    0:temp = 7'b0000000;
    1:temp = 7'b0001010;
    2:temp = 7'b0010100;
    3:temp = 7'b0011110;
    4:temp = 7'b0101000;
    5:temp = 7'b0110010;
    6:temp = 7'b0111100;
    7:temp = 7'b1000110;
    8:temp = 7'b1010000;
    9:temp = 7'b1011010;
endcase
end       

assign ledg = temp + ones;

endmodule 

//сначала забираем десятку у числа
//Смотрим какое число формируют свичи в битках
//от 1 до 9
//Далее мы берем и по прнципу работы BTD добикидываем к ним числа от 0-9
//чтобы сформировать двузначное число
//Далее
//Для примера
//69 = вы снимаем первых четрых свитчей 6, далее по кейсу
//мы закинем 9ку
//Верилог умный, он сам там все преобразует
