module wrap_3 (
    input [7:0] SW,
    output [7:0] LEDG
);

lab_3_3_1 init_1 (SW[7:0], LEDG[7:0]);

endmodule