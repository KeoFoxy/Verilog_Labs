module lab_3_2_1(sw, hex1, y);
input [3:0] sw;
output [6:0] hex1;
output [3:0] y;

wire z;
//Если на свичах больше 9, то на экранчик
//Отвечающий за десятые
//Выводим 1 для чисел 10-19 (1 + число от прошлого задания)
//Если меньше, то пусть остается 0
//И будет срабатывать файл из прошлого задания
//Там уже выводим только 1-9
assign z = (sw[3:0] > 4'b1001);
assign hex1 = (z) ? 7'b1001111 : 7'b1000000;
assign y = (z) ? sw[3:0]-4'b1010 : sw[3:0]; // Забираем единицы из числа
//Надо взять 3 из 13
//Вычтем из 13 10 побитово и почим 3, которую потом запихнем во второй файл
//и там через кейс уже выведем это число в другом файле
//Файлы у нас связаны через оболочку, которая стягивает их
//

endmodule